Joining room 
Går in i rummet 
werewolfbot
varulvsbot
Error when joining room
Kunde inte gå in i rummet
Hi, I am the werewolf bot.
Hej,  jag är varulvsboten.
To join the game, send 'join' to me privately.  List participants with 'who' in public.  To start the game, say 'start' in public.
För att gå med i spelet, skriv 'join' till mig privat.  Få lista på deltagare med 'who' publikt.  För att starta spelet, skriv 'start' publikt.
werewolf
varulv
villager
bybo
 has joined the game.
 har gått med i spelet.
You probably meant 'join'.
Du menade antagligen 'join'.
No players yet.
Inga spelare än.
Not enough players.
Inte tillräckligt med spelare.
You are a werewolf.  
Du är en varulv.  
There are no other werewolves.
Det finns inga andra varulvar.
The other werewolves are: 
De andra varulvarna är: 
You are a villager.
Du är en bybo.
As the sun sets over the little village, the people realize that there is only one side left.  
När solen går ner över den lilla byn, inser folket att det bara finns en sida kvar.  
The villagers have won!
Byborna har vunnit!
The werewolves have won!
Varulvarna har vunnit!
The villagers, tired after the hard work in the fields, go to bed, and the sun sets.  But in the middle of the night, the werewolves wake up!
Byborna, trötta efter dagens hårda arbete, går och lägger sig, och solen går ner.  Men mitt i natten vaknar varulvarna!
You and the other werewolves vote for a villager to kill by typing 'kill NICK' to me.
Du och de andra varulvarna röstar om vilken bybo ni ska döda genom att skriva 'kill NICK' till mig.
A scream of pain and agony is heard!
Ett vrål av smärta och ångest hörs!
 has been devoured by the werewolves.
 har blivit uppäten av varulvarna.
You are not a werewolf.  You are supposed to be sleeping!
Du är ingen varulv.  Du borde sova nu!
 is not a villager.
 är ingen bybo.
 has voted to kill 
 har röstat för att döda 
I don't understand that.
Jag förstår inte.
As the sun rises over the little village, the people realize that there is only one side left.  
När solen går upp över den lilla byn inser folket att det bara finns en sida kvar.
The villagers are outraged over this crime, and want to execute somebody.  They gather in the town square to vote about whom to kill.  Type 'kill NICK' in public to vote.
Byborna är mycket upprörda över detta brott, och vill avrätta någon.  De samlas på torget för att rösta om vem de ska döda.  Skriv 'kill NICK' publikt för att rösta.
The villagers have chosen by simple majority to execute 
Byborna har genom enkelt majoritet valt att avrätta 
All villagers have cast their vote, but no majority has been reached.  The disgruntled villagers go home.
Alla byborna har röstat, men ingen majoritet har uppnåtts.  De missnöjda byborna går hem.
: You are not entitled to vote.
: Du har ingen rösträtt.
 is not a villager.
 är ingen bybo.
